grammar edu:umn:cs:melt:sharedemo:exts:condtable:abstractsyntax;

imports silver:core hiding group;

imports silver:langutil;
imports silver:langutil:pp;

imports edu:umn:cs:melt:sharedemo:host:abstractsyntax;
