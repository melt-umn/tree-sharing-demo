grammar edu:umn:cs:melt:sharedemo:exts:forloop;

exports edu:umn:cs:melt:sharedemo:exts:forloop:concretesyntax;
