grammar edu:umn:cs:melt:sharedemo:host;

imports silver:core;
imports silver:langutil;
imports silver:langutil:pp;
