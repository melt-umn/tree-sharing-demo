grammar edu:umn:cs:melt:sharedemo:translation;

imports silver:core hiding group;

imports edu:umn:cs:melt:sharedemo:host:abstractsyntax;
imports silver:langutil;
imports silver:langutil:pp;
