grammar edu:umn:cs:melt:sharedemo:host;

exports edu:umn:cs:melt:sharedemo:host:concretesyntax;
