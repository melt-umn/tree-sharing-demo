grammar edu:umn:cs:melt:sharedemo:host:abstractsyntax;

imports silver:core;
imports silver:langutil;
imports silver:langutil:pp;
