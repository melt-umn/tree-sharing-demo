grammar edu:umn:cs:melt:sharedemo:exts:condtable;

exports edu:umn:cs:melt:sharedemo:exts:condtable:concretesyntax;
