grammar edu:umn:cs:melt:sharedemo:exts:forloop:abstractsyntax;

imports silver:langutil;
imports silver:langutil:pp;

imports edu:umn:cs:melt:sharedemo:host:abstractsyntax;
imports edu:umn:cs:melt:sharedemo:translation;
